module part1(SW, LEDG);
	input [9:0] SW;
	output [9:0] LEDG;
	
	assign LEDG = SW;
endmodule
